`timescale 1ns / 1ps


module Not(
    input wire a,
    output wire y
    );
    assign y =~a;
endmodule
